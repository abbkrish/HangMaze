module draw_letter #(y=0, x=0, size_y = 20, size_x = 40) (
	input [9:0] DrawX, DrawY,
	input [0:size_x-1] maze_letters [size_y-1:0],
	output draw
	);

	assign draw = ( maze_letters[y][x] && DrawX >= 16*x && (DrawX) < 16*(x+1) && DrawY >= 16*y && DrawY < 16*(y+1) ) ? 1'b1 : 1'b0;
	
endmodule
