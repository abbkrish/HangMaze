module sprite_alphabet (
	input [7:0] sprite_index,
	output [0:15] sprite [15:0]
);

	always_comb
	begin
		unique case (sprite_index)
		8'h00:
		begin
			sprite[0] = 16'b0000000000000000; // 0   yep, this little fucker; he's back
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2 
			sprite[3] = 16'b0000000000000000; // 3 
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000000000000000; // 5
			sprite[6] = 16'b0000000000000000; // 6
			sprite[7] = 16'b0000000000000000; // 7
			sprite[8] = 16'b0000000000000000; // 8
			sprite[9] = 16'b0000000000000000; // 9
			sprite[10] = 16'b0000000000000000; // a
			sprite[11] = 16'b0000000000000000; // b
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000; // f
		end
		8'h01:
		begin
			sprite[0] = 16'b0000000000000000; // 0   yep, this little fucker; he's back
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000011111100000; // 2   ******
			sprite[3] = 16'b0000100000010000; // 3  *      *
			sprite[4] = 16'b0000101001010000; // 4  * *  * *
			sprite[5] = 16'b0000100000010000; // 5  *      *
			sprite[6] = 16'b0000100000010000; // 6  *      *
			sprite[7] = 16'b0000101111010000; // 7  * **** *
			sprite[8] = 16'b0000100110010000; // 8  *  **  *
			sprite[9] = 16'b0000100000010000; // 9  *      *
			sprite[10] = 16'b0000100000010000; // a *      *
			sprite[11] = 16'b0000011111100000; // b  ******
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000; // f
		end
		8'h61:
		begin
			sprite[0] = 16'b0000000000000000; // 0 
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011110000000; // 5  ****
			sprite[6] = 16'b0000000011000000; // 6     **
			sprite[7] = 16'b0000011111000000; // 7  *****
			sprite[8] = 16'b0000110011000000; // 8 **  **
			sprite[9] = 16'b0000110011000000; // 9 **  **
			sprite[10] = 16'b0000110011000000; // a **  **
			sprite[11] = 16'b0000011101100000; // b  *** **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
		
			 // code x62
		8'h62:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000111000000000; // 2  ***
			sprite[3] = 16'b0000011000000000; // 3   **
			sprite[4] = 16'b0000011000000000; // 4   **
			sprite[5] = 16'b0000011110000000; // 5   ****
			sprite[6] = 16'b0000011011000000; // 6   ** **
			sprite[7] = 16'b0000011001100000; // 7   **  **
			sprite[8] = 16'b0000011001100000; // 8   **  **
			sprite[9] = 16'b0000011001100000; // 9   **  **
			sprite[10] = 16'b0000011001100000; // a   **  **
			sprite[11] = 16'b0000011111000000; // b   *****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x63
		8'h63:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011111000000; // 5  *****
			sprite[6] = 16'b0000110001100000; // 6 **   **
			sprite[7] = 16'b0000110000000000; // 7 **
			sprite[8] = 16'b0000110000000000; // 8 **
			sprite[9] = 16'b0000110000000000; // 9 **
			sprite[10] = 16'b0000110001100000; // a **   **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x64
		8'h64:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000111000000; // 2    ***
			sprite[3] = 16'b0000000011000000; // 3     **
			sprite[4] = 16'b0000000011000000; // 4     **
			sprite[5] = 16'b0000001111000000; // 5   ****
			sprite[6] = 16'b0000011011000000; // 6  ** **
			sprite[7] = 16'b0000110011000000; // 7 **  **
			sprite[8] = 16'b0000110011000000; // 8 **  **
			sprite[9] = 16'b0000110011000000; // 9 **  **
			sprite[10] = 16'b0000110011000000; // a **  **
			sprite[11] = 16'b0000011101100000; // b  *** **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x65
		8'h65:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011111000000; // 5  *****
			sprite[6] = 16'b0000110001100000; // 6 **   **
			sprite[7] = 16'b0000111111100000; // 7 *******
			sprite[8] = 16'b0000110000000000; // 8 **
			sprite[9] = 16'b0000110000000000; // 9 **
			sprite[10] = 16'b0000110001100000; // a **   **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x66
		8'h66:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000001110000000; // 2   ***
			sprite[3] = 16'b0000011011000000; // 3  ** **
			sprite[4] = 16'b0000011001000000; // 4  **  *
			sprite[5] = 16'b0000011000000000; // 5  **
			sprite[6] = 16'b0000111100000000; // 6 ****
			sprite[7] = 16'b0000011000000000; // 7  **
			sprite[8] = 16'b0000011000000000; // 8  **
			sprite[9] = 16'b0000011000000000; // 9  **
			sprite[10] = 16'b0000011000000000; // a  **
			sprite[11] = 16'b0000111100000000; // b ****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x67
		8'h67:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011101100000; // 5  *** **
			sprite[6] = 16'b0000110011000000; // 6 **  **
			sprite[7] = 16'b0000110011000000; // 7 **  **
			sprite[8] = 16'b0000110011000000; // 8 **  **
			sprite[9] = 16'b0000110011000000; // 9 **  **
			sprite[10] = 16'b0000110011000000; // a **  **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000000011000000; // c     **
			sprite[13] = 16'b0000110011000000; // d **  **
			sprite[14] = 16'b0000011110000000; // e  ****
			sprite[15] = 16'b0000000000000000;
		end
			 // code x68
		8'h68:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000111000000000; // 2 ***
			sprite[3] = 16'b0000011000000000; // 3  **
			sprite[4] = 16'b0000011000000000; // 4  **
			sprite[5] = 16'b0000011011000000; // 5  ** **
			sprite[6] = 16'b0000011101100000; // 6  *** **
			sprite[7] = 16'b0000011001100000; // 7  **  **
			sprite[8] = 16'b0000011001100000; // 8  **  **
			sprite[9] = 16'b0000011001100000; // 9  **  **
			sprite[10] = 16'b0000011001100000; // a  **  **
			sprite[11] = 16'b0000111001100000; // b ***  **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x69
		8'h69:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000110000000; // 2    **
			sprite[3] = 16'b0000000110000000; // 3    **
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000001110000000; // 5   ***
			sprite[6] = 16'b0000000110000000; // 6    **
			sprite[7] = 16'b0000000110000000; // 7    **
			sprite[8] = 16'b0000000110000000; // 8    **
			sprite[9] = 16'b0000000110000000; // 9    **
			sprite[10] = 16'b0000000110000000; // a    **
			sprite[11] = 16'b0000001111000000; // b   ****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x6a
		8'h6a:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000001100000; // 2      **
			sprite[3] = 16'b0000000001100000; // 3      **
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000000011100000; // 5     ***
			sprite[6] = 16'b0000000001100000; // 6      **
			sprite[7] = 16'b0000000001100000; // 7      **
			sprite[8] = 16'b0000000001100000; // 8      **
			sprite[9] = 16'b0000000001100000; // 9      **
			sprite[10] = 16'b0000000001100000; // a      **
			sprite[11] = 16'b0000000001100000; // b      **
			sprite[12] = 16'b0000011001100000; // c  **  **
			sprite[13] = 16'b0000011001100000; // d  **  **
			sprite[14] = 16'b0000001111000000; // e   ****
			sprite[15] = 16'b0000000000000000;
		end
			 // code x6b0000
		8'h6b:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000111000000000; // 2 ***
			sprite[3] = 16'b0000011000000000; // 3  **
			sprite[4] = 16'b0000011000000000; // 4  **
			sprite[5] = 16'b0000011001100000; // 5  **  **
			sprite[6] = 16'b0000011011000000; // 6  ** **
			sprite[7] = 16'b0000011110000000; // 7  ****
			sprite[8] = 16'b0000011110000000; // 8  ****
			sprite[9] = 16'b0000011011000000; // 9  ** **
			sprite[10] = 16'b0000011001100000; // a  **  **
			sprite[11] = 16'b0000111001100000; // b ***  **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x6c
		8'h6c:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000001110000000; // 2   ***
			sprite[3] = 16'b0000000110000000; // 3    **
			sprite[4] = 16'b0000000110000000; // 4    **
			sprite[5] = 16'b0000000110000000; // 5    **
			sprite[6] = 16'b0000000110000000; // 6    **
			sprite[7] = 16'b0000000110000000; // 7    **
			sprite[8] = 16'b0000000110000000; // 8    **
			sprite[9] = 16'b0000000110000000; // 9    **
			sprite[10] = 16'b0000000110000000; // a    **
			sprite[11] = 16'b0000001111000000; // b   ****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x6d
		8'h6d:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000111001100000; // 5 ***  **
			sprite[6] = 16'b0000111111110000; // 6 ********
			sprite[7] = 16'b0000110110110000; // 7 ** ** **
			sprite[8] = 16'b0000110110110000; // 8 ** ** **
			sprite[9] = 16'b0000110110110000; // 9 ** ** **
			sprite[10] = 16'b0000110110110000; // a ** ** **
			sprite[11] = 16'b0000110110110000; // b ** ** **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x6e
		8'h6e:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110111000000; // 5 ** ***
			sprite[6] = 16'b0000011001100000; // 6  **  **
			sprite[7] = 16'b0000011001100000; // 7  **  **
			sprite[8] = 16'b0000011001100000; // 8  **  **
			sprite[9] = 16'b0000011001100000; // 9  **  **
			sprite[10] = 16'b0000011001100000; // a  **  **
			sprite[11] = 16'b0000011001100000; // b  **  **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x6f
		8'h6f:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011111000000; // 5  *****
			sprite[6] = 16'b0000110001100000; // 6 **   **
			sprite[7] = 16'b0000110001100000; // 7 **   **
			sprite[8] = 16'b0000110001100000; // 8 **   **
			sprite[9] = 16'b0000110001100000; // 9 **   **
			sprite[10] = 16'b0000110001100000; // a **   **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x70
		8'h70:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110111000000; // 5 ** ***
			sprite[6] = 16'b0000011001100000; // 6  **  **
			sprite[7] = 16'b0000011001100000; // 7  **  **
			sprite[8] = 16'b0000011001100000; // 8  **  **
			sprite[9] = 16'b0000011001100000; // 9  **  **
			sprite[10] = 16'b0000011001100000; // a  **  **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000011000000000; // c  **
			sprite[13] = 16'b0000011000000000; // d  **
			sprite[14] = 16'b0000111100000000; // e ****
			sprite[15] = 16'b0000000000000000;
		end
			 // code x71
		8'h71:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011101100000; // 5  *** **
			sprite[6] = 16'b0000110011000000; // 6 **  **
			sprite[7] = 16'b0000110011000000; // 7 **  **
			sprite[8] = 16'b0000110011000000; // 8 **  **
			sprite[9] = 16'b0000110011000000; // 9 **  **
			sprite[10] = 16'b0000110011000000; // a **  **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000000011000000; // c     **
			sprite[13] = 16'b0000000011000000; // d     **
			sprite[14] = 16'b0000000111100000; // e    ****
			sprite[15] = 16'b0000000000000000;
		end
			 // code x72
		8'h72:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110111000000; // 5 ** ***
			sprite[6] = 16'b0000011101100000; // 6  *** **
			sprite[7] = 16'b0000011001100000; // 7  **  **
			sprite[8] = 16'b0000011000000000; // 8  **
			sprite[9] = 16'b0000011000000000; // 9  **
			sprite[10] = 16'b0000011000000000; // a  **
			sprite[11] = 16'b0000111100000000; // b ****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x73
		8'h73:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000011111000000; // 5  *****
			sprite[6] = 16'b0000110001100000; // 6 **   **
			sprite[7] = 16'b0000011000000000; // 7  **
			sprite[8] = 16'b0000001110000000; // 8   ***
			sprite[9] = 16'b0000000011000000; // 9     **
			sprite[10] = 16'b0000110001100000; // a **   **
			sprite[11] = 16'b0000011111000000; // b  *****
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x74
		8'h74:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000100000000; // 2    *
			sprite[3] = 16'b0000001100000000; // 3   **
			sprite[4] = 16'b0000001100000000; // 4   **
			sprite[5] = 16'b0000111111000000; // 5 ******
			sprite[6] = 16'b0000001100000000; // 6   **
			sprite[7] = 16'b0000001100000000; // 7   **
			sprite[8] = 16'b0000001100000000; // 8   **
			sprite[9] = 16'b0000001100000000; // 9   **
			sprite[10] = 16'b0000001101100000; // a   ** **
			sprite[11] = 16'b0000000111000000; // b    ***
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x75
		8'h75:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110011000000; // 5 **  **
			sprite[6] = 16'b0000110011000000; // 6 **  **
			sprite[7] = 16'b0000110011000000; // 7 **  **
			sprite[8] = 16'b0000110011000000; // 8 **  **
			sprite[9] = 16'b0000110011000000; // 9 **  **
			sprite[10] = 16'b0000110011000000; // a **  **
			sprite[11] = 16'b0000011101100000; // b  *** **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x76
		8'h76:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110000110000; // 5 **    **
			sprite[6] = 16'b0000110000110000; // 6 **    **
			sprite[7] = 16'b0000110000110000; // 7 **    **
			sprite[8] = 16'b0000110000110000; // 8 **    **
			sprite[9] = 16'b0000011001100000; // 9  **  **
			sprite[10] = 16'b0000001111000000; // a   ****
			sprite[11] = 16'b0000000110000000; // b    **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x77
		8'h77:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110000110000; // 5 **    **
			sprite[6] = 16'b0000110000110000; // 6 **    **
			sprite[7] = 16'b0000110000110000; // 7 **    **
			sprite[8] = 16'b0000110110110000; // 8 ** ** **
			sprite[9] = 16'b0000110110110000; // 9 ** ** **
			sprite[10] = 16'b0000111111110000; // a ********
			sprite[11] = 16'b0000011001100000; // b  **  **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x78
		8'h78:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110000110000; // 5 **    **
			sprite[6] = 16'b0000011001100000; // 6  **  **
			sprite[7] = 16'b0000001111000000; // 7   ****
			sprite[8] = 16'b0000000110000000; // 8    **
			sprite[9] = 16'b0000001111000000; // 9   ****
			sprite[10] = 16'b0000011001100000; // a  **  **
			sprite[11] = 16'b0000110000110000; // b **    **
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
			 // code x79
		8'h79:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000110001100000; // 5 **   **
			sprite[6] = 16'b0000110001100000; // 6 **   **
			sprite[7] = 16'b0000110001100000; // 7 **   **
			sprite[8] = 16'b0000110001100000; // 8 **   **
			sprite[9] = 16'b0000110001100000; // 9 **   **
			sprite[10] = 16'b0000110001100000; // a **   **
			sprite[11] = 16'b0000011111100000; // b  ******
			sprite[12] = 16'b0000000001100000; // c      **
			sprite[13] = 16'b0000000011000000; // d     **
			sprite[14] = 16'b0000111110000000; // e *****
			sprite[15] = 16'b0000000000000000;
		end
			 // code x7a
		8'h7a:
		begin
			sprite[0] = 16'b0000000000000000; // 0
			sprite[1] = 16'b0000000000000000; // 1
			sprite[2] = 16'b0000000000000000; // 2
			sprite[3] = 16'b0000000000000000; // 3
			sprite[4] = 16'b0000000000000000; // 4
			sprite[5] = 16'b0000111111100000; // 5 *******
			sprite[6] = 16'b0000110011000000; // 6 **  **
			sprite[7] = 16'b0000000110000000; // 7    **
			sprite[8] = 16'b0000001100000000; // 8   **
			sprite[9] = 16'b0000011000000000; // 9  **
			sprite[10] = 16'b0000110001100000; // a **   **
			sprite[11] = 16'b0000111111100000; // b *******
			sprite[12] = 16'b0000000000000000; // c
			sprite[13] = 16'b0000000000000000; // d
			sprite[14] = 16'b0000000000000000; // e
			sprite[15] = 16'b0000000000000000;
		end
		default: 
		begin
			sprite[0] = 16'b0;
			sprite[1] = 16'b0;
			sprite[2] = 16'b0;
			sprite[3] = 16'b0;
			sprite[4] = 16'b0;
			sprite[5] = 16'b0;
			sprite[6] = 16'b0;
			sprite[7] = 16'b0;
			sprite[8] = 16'b0;
			sprite[9] = 16'b0;
			sprite[10] = 16'b0;
			sprite[11] = 16'b0;
			sprite[12] = 16'b0;
			sprite[13] = 16'b0;
			sprite[14] = 16'b0;
			sprite[15] = 16'b0;
		end
	endcase
	
	end
	
endmodule